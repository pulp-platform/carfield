// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Nicole Narr <narrn@student.ethz.ch>
// Christopher Reinwardt <creinwar@student.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Alessandro Ottaviano <aottaviano@iis.ee.ethz.ch>
// Maicol Ciani <maicol.ciano@unibo.it>

// Main testbench for carfield chip. It contains code sequences to boot the
// various islands standalone or in cooperation.

module tb_carfield_chip;

  import uvm_pkg::*;
  import carfield_pkg::*;
  import cheshire_pkg::*;

  carfield_chip_fixture fix();

  // cheshire
  string      chs_preload_elf;
  string      chs_boot_hex;
  string      llc_init_file;
  logic [1:0] boot_mode;
  logic [1:0] preload_mode;
  bit [31:0]  exit_code;
  bit         is_dram;

  // safety island
  string      safed_preload_elf;
  logic       safed_boot_mode;
  bit  [31:0] safed_exit_code;
  bit         safed_exit_status;

  localparam int unsigned SafetyIslandClkEnRegAddr         = 32'h20010070;
  localparam int unsigned SafetyIslandIsolateRegAddr       = 32'h20010040;
  localparam int unsigned SafetyIslandIsolateStatusRegAddr = 32'h20010058;

  // security island
  string      secd_preload_elf;
  string      secd_flash_vmem;
  string      secd_mem_4096;
  string      secd_mem_2048;
  string      secd_mem_512;
  logic       secd_boot_mode;

  // hyperbus
  localparam int unsigned HyperbusTburstMax = 32'h20009008;

  // FP Spatz Cluster
  string      spatzd_preload_elf;
  logic [1:0] spatzd_boot_mode;
  bit  [31:0] spatzd_exit_code;
  bit         spatzd_exit_status;
  doub_bt     spatzd_binary_entry;
  doub_bt     spatzd_reg_value;

  localparam int unsigned SpatzdClkEnRegAddr         = 32'h2001007c;
  localparam int unsigned SpatzdIsolateRegAddr       = 32'h2001004c;
  localparam int unsigned SpatzdIsolateStatusRegAddr = 32'h20010064;

  // pulp cluster
  // Useful register addresses
  localparam int unsigned CarL2StartAddr                      = 32'h7800_0000;
  localparam int unsigned CarDramStartAddr                    = 32'h8000_0000;
  localparam int unsigned PulpdNumCores                       = 12;
  localparam int unsigned PulpdBootAddrL2                     = CarL2StartAddr + 32'h8080;
  localparam int unsigned PulpdBootAddrDram                   = CarDramStartAddr + 32'h8080;
  localparam int unsigned PulpdBootAddr                       = 32'h50200040;
  localparam int unsigned PulpdRetAddr                        = 32'h50200100;
  localparam int unsigned CarSocCtrlPulpdClkEnRegAddr         = 32'h20010078;
  localparam int unsigned CarSocCtrlPulpdIsolateRegAddr       = 32'h20010048;
  localparam int unsigned CarSocCtrlPulpdIsolateStatusRegAddr = 32'h20010060;
  localparam int unsigned CarSocCtrlPulpdFetchEnAddr          = 32'h200100c0;
  localparam int unsigned CarSocCtrlPulpdBootEnAddr           = 32'h200100dc;
  localparam int unsigned CarSocCtrlPulpdBusyAddr             = 32'h200100e4;
  localparam int unsigned CarSocCtrlPulpdEocAddr              = 32'h200100e8;
  // sim variables
  string      pulpd_preload_elf;
  logic [1:0] pulpd_boot_mode;
  bit  [31:0] pulpd_exit_code;
  bit  [31:0] pulpd_ret_val;
  doub_bt     pulpd_binary_entry;
  doub_bt     pulpd_reg_value;

  // MailBox
  parameter logic [31:0] CAR_MBOX_BASE             = 32'h40000000;
  parameter logic [31:0] CAR_NUM_MAILBOXES         = 32'h25;
  parameter logic [31:0] MBOX_INT_SND_STAT_OFFSET  = 32'h00;
  parameter logic [31:0] MBOX_INT_SND_SET_OFFSET   = 32'h04;
  parameter logic [31:0] MBOX_INT_SND_CLR_OFFSET   = 32'h08;
  parameter logic [31:0] MBOX_INT_SND_EN_OFFSET    = 32'h0C;
  parameter logic [31:0] MBOX_INT_RCV_STAT_OFFSET  = 32'h40;
  parameter logic [31:0] MBOX_INT_RCV_SET_OFFSET   = 32'h44;
  parameter logic [31:0] MBOX_INT_RCV_CLR_OFFSET   = 32'h48;
  parameter logic [31:0] MBOX_INT_RCV_EN_OFFSET    = 32'h4C;
  parameter logic [31:0] MBOX_LETTER0_OFFSET       = 32'h80;
  parameter logic [31:0] MBOX_LETTER1_OFFSET       = 32'h84;

  parameter logic [31:0] MBOX_SPATZ_CORE0_ID = 32'h0;
  parameter logic [31:0] MBOX_SPATZ_CORE1_ID = 32'h1;

  parameter int unsigned HyperRstCycles = 120100;

  logic [63:0] unused;

  // bypass pll
  logic       bypass_pll;

  // secure boot mode
  logic       secure_boot;

  // Decide whether to preload hyperram model at time 0
  logic        hyp_user_preload;

  // timing format for $display("...$t..", $realtime)
  initial begin : timing_format
    $timeformat(-9, 0, "ns", 9);
  end : timing_format

  initial begin
    // Fetch plusargs or use safe (fail-fast) defaults
    if (!$value$plusargs("BYPASS_PLL=%d",   bypass_pll))      bypass_pll      = 0;
    if (!$value$plusargs("SECURE_BOOT=%d",  secure_boot))     secure_boot     = 0;
    if (!$value$plusargs("CHS_BOOTMODE=%d", boot_mode))       boot_mode       = 0;
    if (!$value$plusargs("CHS_PRELMODE=%d", preload_mode))    preload_mode    = 0;
    if (!$value$plusargs("CHS_BINARY=%s",   chs_preload_elf)) chs_preload_elf = "";
    if (!$value$plusargs("CHS_IMAGE=%s",    chs_boot_hex))    chs_boot_hex    = "";
    if (!$value$plusargs("LLC_INIT_FILE=%s", llc_init_file))  llc_init_file   = "";

    // PLL bypass
    fix.set_bypass_pll(bypass_pll);

    // Set boot mode and preload boot image if there is one
    fix.set_secure_boot(secure_boot);
    fix.chs_vip.set_boot_mode(boot_mode);
    fix.chs_vip.i2c_eeprom_preload(chs_boot_hex);
    fix.chs_vip.spih_norflash_preload(chs_boot_hex);

    if (chs_preload_elf != "" || chs_boot_hex != "") begin

      // Wait for reset
      fix.chs_vip.wait_for_reset();

    $display("[TB] INFO: Initialize LLC data ways with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[0].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[1].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[2].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[3].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[4].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[5].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[6].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[7].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_0__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_1__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_2__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_3__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_4__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_5__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_6__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_7__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

    $display("[TB] INFO: Initialize L2 memory banks with random values.");
`ifdef CARFIELD_CHIP_NETLIST
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

`ifndef CARFIELD_CHIP_NETLIST
    // initialize the flash info partitions to random values
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[0].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[1].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[2].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[0].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[1].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[2].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[0].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[1].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[2].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[0].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[1].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[2].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
`else
    // initialize the flash info partitions to random values
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_0__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_1__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_2__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_0__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_1__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_2__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_0__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_1__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_2__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_0__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_1__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_2__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
`endif

      // Writing max burst length in Hyperbus configuration registers to
      // prevent the Verification IPs from triggering timing checks.
      $display("[TB] INFO: Configuring Hyperbus through serial link.");
      fix.chs_vip.slink_write_32(HyperbusTburstMax, 32'd128);

      // When Cheshire is offloading to safety island, the latter should be set in passive preloaded
      // bootmode
      fix.safed_vip.set_safed_boot_mode(safety_island_pkg::Preloaded);
      // Preload in idle mode or wait for completion in autonomous boot
      if (boot_mode == 0) begin
        // Idle boot: preload with the specified mode
        case (preload_mode)
          0: begin      // JTAG
            // Cheshire
            is_dram = uvm_re_match("dram",chs_preload_elf);
            if(~is_dram) begin
              $display("Wait the hyperram");
              repeat(HyperRstCycles)
`ifndef CARFIELD_CHIP_NETLIST
                @(posedge fix.i_dut.periph_clk);
`else
                #10ns;
`endif
            end
            fix.chs_vip.jtag_init();
            fix.chs_vip.jtag_elf_run(chs_preload_elf);
            fix.chs_vip.jtag_wait_for_eoc(exit_code);
          end 1: begin  // Standalone Serial Link passive preload
            fix.chs_vip.slink_elf_run(chs_preload_elf);
            fix.chs_vip.slink_wait_for_eoc(exit_code);
          end 2: begin  // Standalone UART passive preload
            fix.chs_vip.uart_debug_elf_run_and_wait(chs_preload_elf, exit_code);
          end 3: begin  // Secure boot: Opentitan booting CVA6
            fix.chs_vip.slink_elf_preload(chs_preload_elf, unused);
            fix.chs_vip.jtag_init();
            fix.chs_vip.jtag_wait_for_eoc(exit_code);
          end default: begin
            $fatal(1, "Unsupported preload mode %d (reserved)!", boot_mode);
          end
        endcase
      end else if (boot_mode == 1) begin
        $fatal(1, "Unsupported boot mode %d (SD Card)!", boot_mode);
      end else begin
        // Autonomous boot: Only poll return code
        fix.chs_vip.jtag_init();
        fix.chs_vip.jtag_wait_for_eoc(exit_code);
      end

      // Sample carfield's clock source frequencies (host, alt, periph)
      //fix.sample_freq_debug_signals();

      // Eventually wait for HWRoT to end initialization and assert Ibex's fetch enable
      fix.passthrough_or_wait_for_secd_hw_init();

      // Wait for the UART to finish reading the current byte
      wait (fix.chs_vip.uart_reading_byte == 0);

      $finish;
    end
  end

  // safety island standalone
  initial begin
    // Fetch plusargs or use safe (fail-fast) defaults
    if (!$value$plusargs("BYPASS_PLL=%d",     bypass_pll))        bypass_pll        = 0;
    if (!$value$plusargs("SECURE_BOOT=%d",    secure_boot))       secure_boot       = 0;
    if (!$value$plusargs("SAFED_BOOTMODE=%d", safed_boot_mode))   safed_boot_mode   = 0;
    if (!$value$plusargs("SAFED_BINARY=%s",   safed_preload_elf)) safed_preload_elf = "";

    // PLL bypass
    fix.set_bypass_pll(bypass_pll);

    // set secure boot mode
    fix.set_secure_boot(secure_boot);

    // set boot mode before reset
    fix.safed_vip.set_safed_boot_mode(safed_boot_mode);

    if (safed_preload_elf != "") begin

      fix.safed_vip.safed_wait_for_reset();

    $display("[TB] INFO: Initialize LLC data ways with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[0].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[1].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[2].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[3].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[4].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[5].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[6].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[7].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_0__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_1__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_2__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_3__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_4__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_5__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_6__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_7__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

    $display("[TB] INFO: Initialize L2 memory banks with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

      // Writing max burst length in Hyperbus configuration registers to
      // prevent the Verification IPs from triggering timing checks.
      $display("[TB] INFO: Configuring Hyperbus through serial link.");
      fix.safed_vip.axi_write_32(HyperbusTburstMax, 32'd128);

      $display("[TB] %t - Enabling safety island clock for stand-alone tests ", $realtime);
      // Clock island after PoR
      fix.safed_vip.axi_write_32(SafetyIslandClkEnRegAddr, 32'h1);
      $display("[TB] %t - De-isolate safety island for stand-alone tests ", $realtime);
      // De-isolate island after PoR
      fix.safed_vip.axi_write_32(SafetyIslandIsolateRegAddr, 32'h0);

      case (safed_boot_mode)
        0: begin
          fix.safed_vip.jtag_safed_init();
          fix.safed_vip.jtag_write_test(32'h6000_1000, 32'hABBA_ABBA);
          fix.safed_vip.jtag_safed_elf_run(safed_preload_elf);
          fix.safed_vip.jtag_safed_wait_for_eoc(safed_exit_code, safed_exit_status);
        end 1: begin
          fix.safed_vip.axi_safed_elf_run(safed_preload_elf);
          fix.safed_vip.axi_safed_wait_for_eoc(safed_exit_code, safed_exit_status);
       end default: begin
          $fatal(1, "Unsupported boot mode %d (reserved)!", safed_boot_mode);
        end
      endcase

      $finish;
    end
  end

  // security island standalone
  initial begin
    // Fetch plusargs or use safe (fail-fast) defaults
    if (!$value$plusargs("BYPASS_PLL=%d",    bypass_pll))       bypass_pll       = 0;
    if (!$value$plusargs("SECURE_BOOT=%d",   secure_boot))      secure_boot      = 0;
    if (!$value$plusargs("SECD_IMAGE=%s",    secd_flash_vmem))  secd_flash_vmem  = "";
    if (!$value$plusargs("SECD_BINARY=%s",   secd_preload_elf)) secd_preload_elf = "";
    if (!$value$plusargs("SECD_MEM_4096=%s", secd_mem_4096 ))   secd_mem_4096    = "";
    if (!$value$plusargs("SECD_MEM_2048=%s", secd_mem_2048 ))   secd_mem_2048    = "";
    if (!$value$plusargs("SECD_MEM_512=%s" , secd_mem_512  ))   secd_mem_512     = "";
    if (!$value$plusargs("SECD_BOOTMODE=%d", secd_boot_mode))   secd_boot_mode   = 0;

    // PLL bypass
    fix.set_bypass_pll(bypass_pll);

    // set secure boot mode
    fix.set_secure_boot(secure_boot);

    // set bootmode
    fix.secd_vip.set_secd_boot_mode(secd_boot_mode);

    if (secd_preload_elf != "" || secd_flash_vmem != "") begin
      // Wait for reset
      fix.chs_vip.wait_for_reset();

    $display("[TB] INFO: Initialize LLC data ways with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[0].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[1].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[2].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[3].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[4].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[5].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[6].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[7].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_0__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_1__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_2__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_3__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_4__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_5__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_6__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_7__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

    $display("[TB] INFO: Initialize L2 memory banks with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

`ifndef CARFIELD_CHIP_NETLIST
    // initialize the flash info partitions to random values
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[0].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[1].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[2].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[0].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[1].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[2].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[0].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[1].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[0].u_prim_flash_bank.gen_info_types[2].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[0].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[1].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.gen_info_types[2].u_info_mem.ram_primitive.gen_2560w_76dw_8be.i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem.i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks[1].u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw.sram_bank_4096w_76dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
`else
    // initialize the flash info partitions to random values
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_0__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_1__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_2__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_0__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_1__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_512,  tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_2__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_512w76b_flash_info_cut.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_512x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_0__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_1__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_0__u_prim_flash_bank.gen_info_types_2__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_0__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_1__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_2048, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.gen_info_types_2__u_info_mem.ram_primitive.gen_2560w_76dw_8be_i_2048w76b_flash_info_cut.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
    $readmemh(secd_mem_4096, tb_carfield_chip.fix.i_dut.i_carfield_soc.gen_secure_subsystem_i_security_island.u_RoT.u_flash_ctrl.u_eflash.u_flash.gen_prim_flash_banks_1__u_prim_flash_bank.u_mem.ram_primitive.gen_32768w_76dw_sram_bank_4096w_76dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x76m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY );
`endif

      // Writing max burst length in Hyperbus configuration registers to
      // prevent the Verification IPs from triggering timing checks.
      $display("[TB] INFO: Configuring Hyperbus through serial link.");
      fix.chs_vip.slink_write_32(HyperbusTburstMax, 32'd128);

      case(secd_boot_mode)
        0: begin
          // Wait before security island HW is initialized
          repeat(10000)
            @(posedge fix.ref_clk);
          fix.secd_vip.debug_secd_module_init();
          fix.secd_vip.load_secd_binary(secd_preload_elf);
          fix.secd_vip.jtag_secd_data_preload();
          fix.secd_vip.jtag_secd_wakeup(32'hE0000080);
          fix.secd_vip.jtag_secd_wait_eoc();
        end 1: begin
          fix.secd_vip.spih_norflash_preload(secd_flash_vmem);
          repeat(10000)
            @(posedge fix.ref_clk);
          fix.secd_vip.jtag_secd_wait_eoc();
        end default: begin
          $fatal(1, "Unsupported boot mode %d (reserved)!", safed_boot_mode);
        end
      endcase
    end
  end

  // pulp cluster standalone
  initial begin
    // Fetch plusargs or use safe (fail-fast) defaults
    if (!$value$plusargs("BYPASS_PLL=%d",         bypass_pll))         bypass_pll        = 0;
    if (!$value$plusargs("PULPD_BOOTMODE=%d",     pulpd_boot_mode))    pulpd_boot_mode   = 0;
    if (!$value$plusargs("PULPD_BINARY=%s",       pulpd_preload_elf))  pulpd_preload_elf = "";
    if (!$value$plusargs("HYP_USER_PRELOAD=%s",   hyp_user_preload))   hyp_user_preload  = 0;

    // PLL bypass
    fix.set_bypass_pll(bypass_pll);

    // Wait for reset
    fix.chs_vip.wait_for_reset();

    if (pulpd_preload_elf != "") begin

    $display("[TB] INFO: Initialize LLC data ways with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[0].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[1].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[2].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[3].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[4].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[5].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[6].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[7].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_0__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_1__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_2__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_3__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_4__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_5__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_6__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_7__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

    $display("[TB] INFO: Initialize L2 memory banks with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

      $display("[TB] %t - Enabling PULP cluster clock for stand-alone tests ", $realtime);
      // Clock island after PoR
      fix.chs_vip.slink_write_32(CarSocCtrlPulpdClkEnRegAddr, 32'h1);
      $display("[TB] %t - De-isolate PULP cluster for stand-alone tests ", $realtime);
      // De-isolate island after PoR
      fix.chs_vip.slink_write_32(CarSocCtrlPulpdIsolateRegAddr, 32'h0);

      case (pulpd_boot_mode)
        0: begin
          // JTAG
          $display("[JTAG PULPD] Init ");
          fix.chs_vip.jtag_init();
          $display("[JTAG PULPD] Halt the core and load the binary to L2 ");
          fix.chs_vip.jtag_elf_halt_load(pulpd_preload_elf, pulpd_binary_entry );

          // boot
          // Write bootaddress to each core
          $display("[JTAG PULPD] Write PULP cluster boot address for each core");
          for (int c = 0; c < PulpdNumCores; c++) begin
            fix.chs_vip.jtag_write_reg32(PulpdBootAddr + c*32'h4, PulpdBootAddrL2);
          end
          // Write boot enable
          $display("[JTAG PULPD] Write PULP cluster boot enable");
          fix.chs_vip.jtag_write_reg32(CarSocCtrlPulpdBootEnAddr, 32'h1);
          // Write fetch enable
          $display("[JTAG PULPD] Write PULP cluster fetch enable");
          fix.chs_vip.jtag_write_reg32(CarSocCtrlPulpdFetchEnAddr, 32'h1);

          // Poll memory address for PULP EOC
          fix.chs_vip.jtag_poll_bit0(CarSocCtrlPulpdEocAddr, pulpd_exit_code, 20);
          fix.slink_read_reg(PulpdRetAddr, pulpd_ret_val, 20);
          if (pulpd_ret_val[30:0] != 'h0) $error("[JTAG PULP] FAILED: return code %x", pulpd_ret_val);
          else $display("[JTAG PULP] SUCCESS");
        end

        1: begin
          // serial link

          // preload
          $display("[SLINK PULPD] Preload the binary to L2 ");
          fix.chs_vip.slink_elf_preload(pulpd_preload_elf, pulpd_binary_entry);

          // boot
          // Write bootaddress to each core
          $display("[SLINK PULPD] Write PULP cluster boot address for each core");
          for (int c = 0; c < PulpdNumCores; c++) begin
            fix.chs_vip.slink_write_32(PulpdBootAddr + c*32'h4, PulpdBootAddrL2);
          end
          // Write boot enable
          $display("[SLINK PULPD] Write PULP cluster boot enable");
          fix.chs_vip.slink_write_32(CarSocCtrlPulpdBootEnAddr, 32'h1);
          // Write fetch enable
          $display("[SLINK PULPD] Write PULP cluster fetch enable");
          fix.chs_vip.slink_write_32(CarSocCtrlPulpdFetchEnAddr, 32'h1);

          // Poll memory address for PULP EOC
          fix.chs_vip.slink_poll_bit0(CarSocCtrlPulpdEocAddr, pulpd_exit_code, 20);
          fix.slink_read_reg(PulpdRetAddr, pulpd_ret_val, 20);
          if (pulpd_ret_val[30:0] != 'h0) $error("[SLINK PULP] FAILED: return code %x", pulpd_ret_val);
          else $display("[SLINK PULP] SUCCESS");
        end
        default: begin
          $fatal(1, "Unsupported boot mode %d (reserved)!", pulpd_boot_mode);
        end
      endcase

      $finish;
    end

    // Fast preload of hyperram
    if (hyp_user_preload != 0 && pulpd_preload_elf == "") begin
      $warning( "[TB] - Instantly preload hyperram0 and hyperrram1 models at time 0. This preload \
                mode should be used for simulation only, because it does not check whether we can \
                preload the hyperram using physical interfaces, e.g., JTAG or SL. If there is enough \
                confidence physical interfaces are working correctly with a gate-level netlist, this \
                mode could be used to speed up the simulation, but at your own risk. You were \
                warned. \n");
      // Hyperrams models are preloaded at time 0. Preferably, this bootflow is used with cluster
      // accelerators, but can be extended to other islands as well. We check the EOC with the JTAG

      $display("[TB] %t - Wait for HyperRAM", $realtime);
      repeat(HyperRstCycles)
`ifndef CARFIELD_CHIP_NETLIST
        @(posedge fix.i_dut.periph_clk);
`else
        #10ns;
`endif

      $display("[TB] %t - Enabling PULP cluster clock for stand-alone tests ", $realtime);
      // Clock island after PoR
      fix.chs_vip.slink_write_32(CarSocCtrlPulpdClkEnRegAddr, 32'h1);
      $display("[TB] %t - De-isolate PULP cluster for stand-alone tests ", $realtime);
      // De-isolate island after PoR
      fix.chs_vip.slink_write_32(CarSocCtrlPulpdIsolateRegAddr, 32'h0);

      // Write bootaddress to each core
      $display("[SLINK PULPD] Write PULP cluster boot address for each core");
      for (int c = 0; c < PulpdNumCores; c++) begin
        fix.chs_vip.slink_write_32(PulpdBootAddr + c*32'h4, PulpdBootAddrDram);
      end
      // Write boot enable
      $display("[SLINK PULPD] Write PULP cluster boot enable");
      fix.chs_vip.slink_write_32(CarSocCtrlPulpdBootEnAddr, 32'h1);
      // Write fetch enable
      $display("[SLINK PULPD] Write PULP cluster fetch enable");
      fix.chs_vip.slink_write_32(CarSocCtrlPulpdFetchEnAddr, 32'h1);

      // Poll memory address for PULP EOC
      fix.chs_vip.slink_poll_bit0(CarSocCtrlPulpdEocAddr, pulpd_exit_code, 20);
      fix.slink_read_reg(PulpdRetAddr, pulpd_ret_val, 20);
      if (pulpd_ret_val[30:0] != 'h0) $error("[JTAG PULP] FAILED: return code %x", pulpd_ret_val);
      else $display("[SLINK PULP] SUCCESS");

      $finish;
    end
  end

  // spatz cluster standalone
  initial begin
    // Fetch plusargs or use safe (fail-fast) defaults
    if (!$value$plusargs("BYPASS_PLL=%d",     bypass_pll))        bypass_pll        = 0;
    if (!$value$plusargs("SECURE_BOOT=%d",     secure_boot))        secure_boot        = 0;
    if (!$value$plusargs("SPATZD_BOOTMODE=%d", spatzd_boot_mode))   spatzd_boot_mode   = 0;
    if (!$value$plusargs("SPATZD_BINARY=%s",   spatzd_preload_elf)) spatzd_preload_elf = "";

    // PLL bypass
    fix.set_bypass_pll(bypass_pll);

    // set secure boot mode
    fix.set_secure_boot(secure_boot);

    if (spatzd_preload_elf != "") begin

      // Wait for reset
      fix.chs_vip.wait_for_reset();

    $display("[TB] INFO: Initialize LLC data ways with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[0].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[1].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[2].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[3].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[4].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[5].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[6].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc.i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways[7].i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be.sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_0__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_1__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_2__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_3__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_4__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_5__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_6__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh(llc_init_file, tb_carfield_chip.fix.i_dut.i_carfield_soc.i_cheshire_wrap.i_cheshire_soc.gen_llc_i_llc.i_axi_llc_top_raw.i_llc_ways.gen_data_ways_7__i_data_way.i_data_sram.i_data_sram.gen_2048w_64dw_8be_sram_bank_2048w_64dw.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_2048x64m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

    $display("[TB] INFO: Initialize L2 memory banks with random values.");
`ifndef CARFIELD_CHIP_NETLIST
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[0].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[0].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[0].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[1].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[2].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[3].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[4].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[5].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[6].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[7].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[8].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[9].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[10].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[11].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[12].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[13].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[14].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group[1].i_car_l2_bank_group.genblk1[1].i_ecc_sram_wrap.i_bank.gen_65536w_39dw.sram_bank_4096w_39dw_cut[15].i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`else
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_0__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_0__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);

      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_0__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_1__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_2__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_3__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_4__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_5__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_6__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_7__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_8__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_9__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_10__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_11__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_12__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_13__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_14__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
      $readmemh("/usr/scratch2/fenga9/lbertaccini/carfield-pd-mr/l2_init_file.vmem", tb_carfield_chip.fix.i_dut.i_carfield_soc.i_reconfigurable_l2.i_l2_top.gen_bank_group_1__i_car_l2_bank_group.genblk1_1__i_ecc_sram_wrap.i_bank.gen_65536w_39dw_sram_bank_4096w_39dw_cut_15__i_cut.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_bmod.ip224uhdlp1p11rf_4096x39m4b2c1s1_t0r0p0d0a1m1h_array.DATA_ARRAY);
`endif

      // Writing max burst length in Hyperbus configuration registers to
      // prevent the Verification IPs from triggering timing checks.
      $display("[TB] INFO: Configuring Hyperbus through serial link.");
      fix.chs_vip.slink_write_32(HyperbusTburstMax, 32'd128);

      $display("[TB] %t - Enabling spatz clock for stand-alone tests ", $realtime);
      // Clock island after PoR
      fix.chs_vip.slink_write_32(SpatzdClkEnRegAddr, 32'h1);
      $display("[TB] %t - De-isolate spatz for stand-alone tests ", $realtime);
      // De-isolate island after PoR
      fix.chs_vip.slink_write_32(SpatzdIsolateRegAddr, 32'h0);

      case (spatzd_boot_mode)
        0: begin
          // JTAG
          $display("[JTAG SPATZD] Init ");
          fix.chs_vip.jtag_init();
          $display("[JTAG SPATZD] Halt the core and load the binary to L2 ");
          fix.chs_vip.jtag_elf_halt_load(spatzd_preload_elf, spatzd_binary_entry );

          // write start address into the csr
          $display("[JTAG SPATZD] write the CSR %x of spatz with the entry point %x", spatz_cluster_pkg::PeriStartAddr + spatz_cluster_peripheral_reg_pkg::SPATZ_CLUSTER_PERIPHERAL_CLUSTER_BOOT_CONTROL_OFFSET, spatzd_binary_entry);
          fix.chs_vip.jtag_write_reg(spatz_cluster_pkg::PeriStartAddr + spatz_cluster_peripheral_reg_pkg::SPATZ_CLUSTER_PERIPHERAL_CLUSTER_BOOT_CONTROL_OFFSET, spatzd_binary_entry );

          // Set interrupt on mailbox mailbox id MBOX_SPATZD_CORE0_ID and MBOX_SPATZD_CORE1_ID
          spatzd_reg_value = 64'h1;
          $display("[JTAG SPATZD] Set mailbox interrupt ID  %x at %x ",MBOX_SPATZ_CORE0_ID, CAR_MBOX_BASE +  MBOX_INT_SND_SET_OFFSET + (MBOX_SPATZ_CORE0_ID*32'h100));
          fix.chs_vip.jtag_write_reg32(CAR_MBOX_BASE +  MBOX_INT_SND_SET_OFFSET + (MBOX_SPATZ_CORE0_ID*32'h100) , spatzd_reg_value);

          $display("[JTAG SPATZD] Set mailbox interrupt ID  %x at %x ",MBOX_SPATZ_CORE1_ID, CAR_MBOX_BASE +  MBOX_INT_SND_SET_OFFSET + (MBOX_SPATZ_CORE1_ID*32'h100));
          fix.chs_vip.jtag_write_reg32(CAR_MBOX_BASE +  MBOX_INT_SND_SET_OFFSET + (MBOX_SPATZ_CORE1_ID*32'h100) , spatzd_reg_value);

          // Enable interrupt on mailbox id MBOX_SPATZ_CORE0_ID and MBOX_SPATZ_CORE1_ID
          $display("[JTAG SPATZD] Enable mailbox interrupt ID  %x at %x ",MBOX_SPATZ_CORE0_ID, CAR_MBOX_BASE +  MBOX_INT_SND_EN_OFFSET + (MBOX_SPATZ_CORE0_ID*32'h100) ,spatzd_reg_value);
          fix.chs_vip.jtag_write_reg32(CAR_MBOX_BASE +  MBOX_INT_SND_EN_OFFSET + (MBOX_SPATZ_CORE0_ID*32'h100) , spatzd_reg_value);

          $display("[JTAG SPATZD] Enable mailbox interrupt ID  %x at %x ",MBOX_SPATZ_CORE1_ID, CAR_MBOX_BASE +  MBOX_INT_SND_EN_OFFSET + (MBOX_SPATZ_CORE1_ID*32'h100) ,spatzd_reg_value);
          fix.chs_vip.jtag_write_reg32(CAR_MBOX_BASE +  MBOX_INT_SND_EN_OFFSET + (MBOX_SPATZ_CORE1_ID*32'h100) , spatzd_reg_value);

          // Poll memory address for Spatz EOC
          fix.chs_vip.jtag_poll_bit0(spatz_cluster_pkg::PeriStartAddr + spatz_cluster_peripheral_reg_pkg::SPATZ_CLUSTER_PERIPHERAL_CLUSTER_EOC_EXIT_OFFSET, spatzd_exit_code, 20);
          spatzd_exit_code >>= 1;
          if (spatzd_exit_code) $error("[JTAG SPATZ] FAILED: return code %0d", spatzd_exit_code);
          else $display("[JTAG SPATZD] SUCCESS");
        end

        1: begin
          // SERIAL LINK
          $display("[SLINK SPATZD] Preload the binary to L2 ");
          fix.chs_vip.slink_elf_preload(spatzd_preload_elf, spatzd_binary_entry);

          // write start address into the csr
          $display("[SLINK SPATZD] Write the CSR %x of spatz with the entry point %x", spatz_cluster_pkg::PeriStartAddr + spatz_cluster_peripheral_reg_pkg::SPATZ_CLUSTER_PERIPHERAL_CLUSTER_BOOT_CONTROL_OFFSET, spatzd_binary_entry);
          fix.chs_vip.slink_write_32(spatz_cluster_pkg::PeriStartAddr + spatz_cluster_peripheral_reg_pkg::SPATZ_CLUSTER_PERIPHERAL_CLUSTER_BOOT_CONTROL_OFFSET, spatzd_binary_entry);

          // Set interrupt on mailbox ids MBOX_SPATZ_CORE0_ID and MBOX_SPATZ_CORE1_ID
          spatzd_reg_value = 64'h1;
          $display("[SLINK SPATZD] Set mailbox interrupt ID  %x at %x ",MBOX_SPATZ_CORE0_ID, CAR_MBOX_BASE +  MBOX_INT_SND_SET_OFFSET + (MBOX_SPATZ_CORE0_ID*32'h100));
          fix.chs_vip.slink_write_32(CAR_MBOX_BASE +  MBOX_INT_SND_SET_OFFSET + (MBOX_SPATZ_CORE0_ID*32'h100) , spatzd_reg_value);

          $display("[SLINK SPATZD] Set mailbox interrupt ID  %x at %x ",MBOX_SPATZ_CORE0_ID, CAR_MBOX_BASE +  MBOX_INT_SND_SET_OFFSET + (MBOX_SPATZ_CORE1_ID*32'h100));
          fix.chs_vip.slink_write_32(CAR_MBOX_BASE +  MBOX_INT_SND_SET_OFFSET + (MBOX_SPATZ_CORE1_ID*32'h100) , spatzd_reg_value);

          // Enable interrupt on mailbox ids MBOX_SPATZ_CORE0_ID and MBOX_SPATZ_CORE1_ID
          $display("[SLINK SPATZD] Enable mailbox interrupt ID  %x at %x ",MBOX_SPATZ_CORE0_ID, CAR_MBOX_BASE +  MBOX_INT_SND_EN_OFFSET + (MBOX_SPATZ_CORE0_ID*32'h100) ,spatzd_reg_value);
          fix.chs_vip.slink_write_32(CAR_MBOX_BASE +  MBOX_INT_SND_EN_OFFSET + (MBOX_SPATZ_CORE0_ID*32'h100) , spatzd_reg_value);

          $display("[SLINK SPATZD] Enable mailbox interrupt ID  %x at %x ",MBOX_SPATZ_CORE0_ID, CAR_MBOX_BASE +  MBOX_INT_SND_EN_OFFSET + (MBOX_SPATZ_CORE1_ID*32'h100) ,spatzd_reg_value);
          fix.chs_vip.slink_write_32(CAR_MBOX_BASE +  MBOX_INT_SND_EN_OFFSET + (MBOX_SPATZ_CORE1_ID*32'h100) , spatzd_reg_value);

          // Poll memory address for Spatz EOC
          fix.chs_vip.slink_poll_bit0(spatz_cluster_pkg::PeriStartAddr + spatz_cluster_peripheral_reg_pkg::SPATZ_CLUSTER_PERIPHERAL_CLUSTER_EOC_EXIT_OFFSET, spatzd_exit_code, 20);
          spatzd_exit_code >>= 1;
          if (spatzd_exit_code) $error("[SLINK SPATZ] FAILED: return code %0d", spatzd_exit_code);
          else $display("[SLINK SPATZ] SUCCESS");
        end

        default: begin
          $fatal(1, "Unsupported boot mode %d (reserved)!", spatzd_boot_mode);
        end
      endcase
      $finish;
    end
  end

endmodule

